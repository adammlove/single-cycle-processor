module adder_tb(a, b, cin, cout, sum);
  output reg [63:0] a, b;
  output reg cin;
  input wire cout;
  input wire overflow;
  output wire [63:0] sum;
  
  reg [63:0] sum_expected;
  reg cout_expected;
  reg overflow_expected;
  
  reg [31:0] vectornum, errors;
  reg [194:0] testvectors[10000:0];
  
  reg clk, reset;
  
  // initialize the module
  sixtyfourbitadder adder(a, b, cin, cout, overflow, sum);
  
  // generate a clock signal
  always begin
    clk = 0; #5; clk = 1; #5;
  end
  
  // read in a test vector
  initial begin
    $readmemb("adder_testvectors.tv", testvectors);
  	vectornum = 0; errors = 0;
  	reset = 1; #27; reset = 0;
  end
  
  // assign test values
  always @(posedge clk) begin
    #1; {a, b, cin, cout_expected, sum_expected} <= testvectors[vectornum];
  end
  
  // test the values
  always @(negedge clk) begin
    if(~reset)
      begin
        // check the values generated by the module against golden values
        if(sum != sum_expected || cout != cout_expected)
        begin
          $display("%b + %b + %b = %b %b != %b %b", cin, a, b, cout_expected, sum_expected, cout, sum);
          errors <= errors + 1;
        end
        vectornum <= vectornum + 1;

        // once all vectors have been checked
        if(testvectors[vectornum] === 194'bx)
          begin
            $display("finished with %0d errors", errors);
            $finish;
          end
      end
  end
endmodule